module iopll (
		input  wire  refclk,   //  refclk.clk
		output wire  locked,   //  locked.export
		input  wire  rst,      //   reset.reset
		output wire  outclk_0, // outclk0.clk
		output wire  outclk_1  // outclk1.clk
	);
endmodule

