module q_sys_systemclk_f_0 (
		output wire  out_systempll_synthlock_0, // out_systempll_synthlock_0.out_systempll_synthlock
		output wire  out_systempll_clk_0,       //       out_systempll_clk_0.clk
		output wire  out_refclk_fgt_4,          //          out_refclk_fgt_4.clk
		input  wire  in_refclk_fgt_4,           //                refclk_fgt.in_refclk_fgt_4
		input  wire  disable_refclk_monitor_4   //  disable_refclk_monitor_4.disable_refclk_monitor_4
	);
endmodule

